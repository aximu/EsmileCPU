`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/01/01 10:27:51
// Design Name: 
// Module Name: esmilecpu_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "../core/define.v"

module esmilecpu_top(

    input wire  clk,
    input wire  rstn,

    input wire
    input wire 
    input wire 
    input wire 
    input wire 
    input wire 
    input wire 
    input wire 
    input wire 
    );
endmodule
